module grayCode
  (
   input wire[3:0] in,
   output wire[3:0] gray
   );

   assign gray = (in==4'b0000) ? 4'b0000 :
		 (in==4'b0001) ? 4'b0001 :
		 (in==4'b0010) ? 4'b0011 :
		 (in==4'b0011) ? 4'b0010 :
		 (in==4'b0100) ? 4'b0110 :
		 (in==4'b0101) ? 4'b0111 :
		 (in==4'b0110) ? 4'b0101 :
		 (in==4'b0111) ? 4'b0100 :
		 (in==4'b1000) ? 4'b1100 :
		 (in==4'b1001) ? 4'b1101 :
		 (in==4'b1010) ? 4'b1111 :
		 (in==4'b1011) ? 4'b1110 :
		 (in==4'b1100) ? 4'b1010 :
		 (in==4'b1101) ? 4'b1011 :
		 (in==4'b1110) ? 4'b1001 :
		 4'b1000;
endmodule
